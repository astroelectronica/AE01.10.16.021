.title KiCad schematic
.include "models/BSS138W.spice.txt"
.include "models/C2012X7R2A104K125AA_p.mod"
.include "models/CGA4C2C0G1H103J060AD_p.mod"
.include "models/MMBD4148.spice.txt"
.include "models/TLC2272.LIB"
R1 VDD /NTC {Rntc}
R2 /NTC 0 13k
R3 VDD /HYST2V65 20k
R4 /HYST2V65 /TEMP 8.06k
R5 /TEMP 0 11.8k
R6 VDD /HYST0V1 33.2k
R7 /HYST0V1 0 20k
V1 VDD 0 5
XU2 /TRI /HYST0V1 VDD 0 /HYST TLC2272
R8 /HYST0V1 /DRAIN 1.62k
R10 /INTEG /HYST 274k
XU6 /HYST2V65 /INTEG VDD 0 /TRI TLC2272
XU5 /TRI /INTEG CGA4C2C0G1H103J060AD_p
XU7 /COMP /TRI VDD 0 /OUT TLC2272
R9 /K /NTC 3.83k
XU4 /COMP 0 CGA4C2C0G1H103J060AD_p
R11 /COMP 0 40.2k
R12 /CTRL /COMP 162k
V2 /CTRL 0 {VDIMM}
R13 /OUT 0 10k
XU1 /DRAIN /HYST 0 BSS138W
XU3 /TEMP /NTC VDD 0 /K TLC2272
D1 /COMP /K DI_MMBD4148
XU8 VDD 0 C2012X7R2A104K125AA_p
XU9 VDD 0 C2012X7R2A104K125AA_p
.end
